module stream_idct (
      nasti_stream_channel.slave  in_ch,
      nasti_stream_channel.master out_ch,

      input aclk,
      input aresetn
   );

   localparam COEF_WIDTH = 16;

   // In/Out staging registers.
   logic signed [COEF_WIDTH - 1:0] row_idct_in    [0:7];
   logic signed [COEF_WIDTH + 3:0] row_idct_out   [0:7];
   logic signed [COEF_WIDTH - 1:0] row_idct_out_h [0:7];
   logic idct_en, lock_idct, busy_idct, out_en;

   // This is used to perform signed truncation to avoid array size mismatches.
   assign row_idct_out_h[0] = row_idct_out[0];
   assign row_idct_out_h[1] = row_idct_out[1];
   assign row_idct_out_h[2] = row_idct_out[2];
   assign row_idct_out_h[3] = row_idct_out[3];
   assign row_idct_out_h[4] = row_idct_out[4];
   assign row_idct_out_h[5] = row_idct_out[5];
   assign row_idct_out_h[6] = row_idct_out[6];
   assign row_idct_out_h[7] = row_idct_out[7];

   stream_dct_handler handler(
      .in_ch(in_ch),
      .out_ch(out_ch),

      .row_dct_in(row_idct_in),
      .row_dct_out(row_idct_out_h),
      .dct_en(idct_en),
      .lock_dct(lock_idct),
      .busy_dct(busy_idct),
      .out_en(out_en),

      .aclk(aclk),
      .aresetn(aresetn)
   );

   // IDCT Pipeline
   pipelined_idct #(
      .COEF_WIDTH(COEF_WIDTH)
   ) idct_pl(
      .row(row_idct_in),
      .idct_row(row_idct_out),

      .en(idct_en),
      .aclk(aclk),
      .aresetn(aresetn),
      .locked(lock_idct),
      .busy(busy_idct),
      .out_en(out_en)
   );
endmodule
